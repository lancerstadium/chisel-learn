module FileReader(
  input        clock,
  input        reset,
  input  [7:0] io_addr,
  output [7:0] io_data
);
  wire [7:0] _GEN_1 = 8'h1 == io_addr ? 8'h3 : 8'h1; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_2 = 8'h2 == io_addr ? 8'h5 : _GEN_1; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_3 = 8'h3 == io_addr ? 8'h7 : _GEN_2; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_4 = 8'h4 == io_addr ? 8'h9 : _GEN_3; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_5 = 8'h5 == io_addr ? 8'hb : _GEN_4; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_6 = 8'h6 == io_addr ? 8'hd : _GEN_5; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_7 = 8'h7 == io_addr ? 8'hf : _GEN_6; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_8 = 8'h8 == io_addr ? 8'h0 : _GEN_7; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_9 = 8'h9 == io_addr ? 8'h0 : _GEN_8; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_10 = 8'ha == io_addr ? 8'h0 : _GEN_9; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_11 = 8'hb == io_addr ? 8'h0 : _GEN_10; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_12 = 8'hc == io_addr ? 8'h0 : _GEN_11; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_13 = 8'hd == io_addr ? 8'h0 : _GEN_12; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_14 = 8'he == io_addr ? 8'h0 : _GEN_13; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_15 = 8'hf == io_addr ? 8'h0 : _GEN_14; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_16 = 8'h10 == io_addr ? 8'h0 : _GEN_15; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_17 = 8'h11 == io_addr ? 8'h0 : _GEN_16; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_18 = 8'h12 == io_addr ? 8'h0 : _GEN_17; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_19 = 8'h13 == io_addr ? 8'h0 : _GEN_18; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_20 = 8'h14 == io_addr ? 8'h0 : _GEN_19; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_21 = 8'h15 == io_addr ? 8'h0 : _GEN_20; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_22 = 8'h16 == io_addr ? 8'h0 : _GEN_21; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_23 = 8'h17 == io_addr ? 8'h0 : _GEN_22; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_24 = 8'h18 == io_addr ? 8'h0 : _GEN_23; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_25 = 8'h19 == io_addr ? 8'h0 : _GEN_24; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_26 = 8'h1a == io_addr ? 8'h0 : _GEN_25; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_27 = 8'h1b == io_addr ? 8'h0 : _GEN_26; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_28 = 8'h1c == io_addr ? 8'h0 : _GEN_27; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_29 = 8'h1d == io_addr ? 8'h0 : _GEN_28; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_30 = 8'h1e == io_addr ? 8'h0 : _GEN_29; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_31 = 8'h1f == io_addr ? 8'h0 : _GEN_30; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_32 = 8'h20 == io_addr ? 8'h0 : _GEN_31; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_33 = 8'h21 == io_addr ? 8'h0 : _GEN_32; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_34 = 8'h22 == io_addr ? 8'h0 : _GEN_33; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_35 = 8'h23 == io_addr ? 8'h0 : _GEN_34; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_36 = 8'h24 == io_addr ? 8'h0 : _GEN_35; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_37 = 8'h25 == io_addr ? 8'h0 : _GEN_36; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_38 = 8'h26 == io_addr ? 8'h0 : _GEN_37; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_39 = 8'h27 == io_addr ? 8'h0 : _GEN_38; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_40 = 8'h28 == io_addr ? 8'h0 : _GEN_39; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_41 = 8'h29 == io_addr ? 8'h0 : _GEN_40; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_42 = 8'h2a == io_addr ? 8'h0 : _GEN_41; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_43 = 8'h2b == io_addr ? 8'h0 : _GEN_42; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_44 = 8'h2c == io_addr ? 8'h0 : _GEN_43; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_45 = 8'h2d == io_addr ? 8'h0 : _GEN_44; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_46 = 8'h2e == io_addr ? 8'h0 : _GEN_45; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_47 = 8'h2f == io_addr ? 8'h0 : _GEN_46; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_48 = 8'h30 == io_addr ? 8'h0 : _GEN_47; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_49 = 8'h31 == io_addr ? 8'h0 : _GEN_48; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_50 = 8'h32 == io_addr ? 8'h0 : _GEN_49; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_51 = 8'h33 == io_addr ? 8'h0 : _GEN_50; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_52 = 8'h34 == io_addr ? 8'h0 : _GEN_51; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_53 = 8'h35 == io_addr ? 8'h0 : _GEN_52; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_54 = 8'h36 == io_addr ? 8'h0 : _GEN_53; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_55 = 8'h37 == io_addr ? 8'h0 : _GEN_54; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_56 = 8'h38 == io_addr ? 8'h0 : _GEN_55; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_57 = 8'h39 == io_addr ? 8'h0 : _GEN_56; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_58 = 8'h3a == io_addr ? 8'h0 : _GEN_57; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_59 = 8'h3b == io_addr ? 8'h0 : _GEN_58; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_60 = 8'h3c == io_addr ? 8'h0 : _GEN_59; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_61 = 8'h3d == io_addr ? 8'h0 : _GEN_60; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_62 = 8'h3e == io_addr ? 8'h0 : _GEN_61; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_63 = 8'h3f == io_addr ? 8'h0 : _GEN_62; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_64 = 8'h40 == io_addr ? 8'h0 : _GEN_63; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_65 = 8'h41 == io_addr ? 8'h0 : _GEN_64; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_66 = 8'h42 == io_addr ? 8'h0 : _GEN_65; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_67 = 8'h43 == io_addr ? 8'h0 : _GEN_66; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_68 = 8'h44 == io_addr ? 8'h0 : _GEN_67; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_69 = 8'h45 == io_addr ? 8'h0 : _GEN_68; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_70 = 8'h46 == io_addr ? 8'h0 : _GEN_69; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_71 = 8'h47 == io_addr ? 8'h0 : _GEN_70; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_72 = 8'h48 == io_addr ? 8'h0 : _GEN_71; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_73 = 8'h49 == io_addr ? 8'h0 : _GEN_72; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_74 = 8'h4a == io_addr ? 8'h0 : _GEN_73; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_75 = 8'h4b == io_addr ? 8'h0 : _GEN_74; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_76 = 8'h4c == io_addr ? 8'h0 : _GEN_75; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_77 = 8'h4d == io_addr ? 8'h0 : _GEN_76; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_78 = 8'h4e == io_addr ? 8'h0 : _GEN_77; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_79 = 8'h4f == io_addr ? 8'h0 : _GEN_78; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_80 = 8'h50 == io_addr ? 8'h0 : _GEN_79; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_81 = 8'h51 == io_addr ? 8'h0 : _GEN_80; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_82 = 8'h52 == io_addr ? 8'h0 : _GEN_81; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_83 = 8'h53 == io_addr ? 8'h0 : _GEN_82; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_84 = 8'h54 == io_addr ? 8'h0 : _GEN_83; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_85 = 8'h55 == io_addr ? 8'h0 : _GEN_84; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_86 = 8'h56 == io_addr ? 8'h0 : _GEN_85; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_87 = 8'h57 == io_addr ? 8'h0 : _GEN_86; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_88 = 8'h58 == io_addr ? 8'h0 : _GEN_87; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_89 = 8'h59 == io_addr ? 8'h0 : _GEN_88; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_90 = 8'h5a == io_addr ? 8'h0 : _GEN_89; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_91 = 8'h5b == io_addr ? 8'h0 : _GEN_90; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_92 = 8'h5c == io_addr ? 8'h0 : _GEN_91; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_93 = 8'h5d == io_addr ? 8'h0 : _GEN_92; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_94 = 8'h5e == io_addr ? 8'h0 : _GEN_93; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_95 = 8'h5f == io_addr ? 8'h0 : _GEN_94; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_96 = 8'h60 == io_addr ? 8'h0 : _GEN_95; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_97 = 8'h61 == io_addr ? 8'h0 : _GEN_96; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_98 = 8'h62 == io_addr ? 8'h0 : _GEN_97; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_99 = 8'h63 == io_addr ? 8'h0 : _GEN_98; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_100 = 8'h64 == io_addr ? 8'h0 : _GEN_99; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_101 = 8'h65 == io_addr ? 8'h0 : _GEN_100; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_102 = 8'h66 == io_addr ? 8'h0 : _GEN_101; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_103 = 8'h67 == io_addr ? 8'h0 : _GEN_102; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_104 = 8'h68 == io_addr ? 8'h0 : _GEN_103; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_105 = 8'h69 == io_addr ? 8'h0 : _GEN_104; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_106 = 8'h6a == io_addr ? 8'h0 : _GEN_105; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_107 = 8'h6b == io_addr ? 8'h0 : _GEN_106; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_108 = 8'h6c == io_addr ? 8'h0 : _GEN_107; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_109 = 8'h6d == io_addr ? 8'h0 : _GEN_108; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_110 = 8'h6e == io_addr ? 8'h0 : _GEN_109; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_111 = 8'h6f == io_addr ? 8'h0 : _GEN_110; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_112 = 8'h70 == io_addr ? 8'h0 : _GEN_111; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_113 = 8'h71 == io_addr ? 8'h0 : _GEN_112; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_114 = 8'h72 == io_addr ? 8'h0 : _GEN_113; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_115 = 8'h73 == io_addr ? 8'h0 : _GEN_114; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_116 = 8'h74 == io_addr ? 8'h0 : _GEN_115; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_117 = 8'h75 == io_addr ? 8'h0 : _GEN_116; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_118 = 8'h76 == io_addr ? 8'h0 : _GEN_117; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_119 = 8'h77 == io_addr ? 8'h0 : _GEN_118; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_120 = 8'h78 == io_addr ? 8'h0 : _GEN_119; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_121 = 8'h79 == io_addr ? 8'h0 : _GEN_120; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_122 = 8'h7a == io_addr ? 8'h0 : _GEN_121; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_123 = 8'h7b == io_addr ? 8'h0 : _GEN_122; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_124 = 8'h7c == io_addr ? 8'h0 : _GEN_123; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_125 = 8'h7d == io_addr ? 8'h0 : _GEN_124; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_126 = 8'h7e == io_addr ? 8'h0 : _GEN_125; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_127 = 8'h7f == io_addr ? 8'h0 : _GEN_126; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_128 = 8'h80 == io_addr ? 8'h0 : _GEN_127; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_129 = 8'h81 == io_addr ? 8'h0 : _GEN_128; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_130 = 8'h82 == io_addr ? 8'h0 : _GEN_129; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_131 = 8'h83 == io_addr ? 8'h0 : _GEN_130; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_132 = 8'h84 == io_addr ? 8'h0 : _GEN_131; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_133 = 8'h85 == io_addr ? 8'h0 : _GEN_132; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_134 = 8'h86 == io_addr ? 8'h0 : _GEN_133; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_135 = 8'h87 == io_addr ? 8'h0 : _GEN_134; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_136 = 8'h88 == io_addr ? 8'h0 : _GEN_135; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_137 = 8'h89 == io_addr ? 8'h0 : _GEN_136; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_138 = 8'h8a == io_addr ? 8'h0 : _GEN_137; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_139 = 8'h8b == io_addr ? 8'h0 : _GEN_138; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_140 = 8'h8c == io_addr ? 8'h0 : _GEN_139; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_141 = 8'h8d == io_addr ? 8'h0 : _GEN_140; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_142 = 8'h8e == io_addr ? 8'h0 : _GEN_141; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_143 = 8'h8f == io_addr ? 8'h0 : _GEN_142; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_144 = 8'h90 == io_addr ? 8'h0 : _GEN_143; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_145 = 8'h91 == io_addr ? 8'h0 : _GEN_144; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_146 = 8'h92 == io_addr ? 8'h0 : _GEN_145; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_147 = 8'h93 == io_addr ? 8'h0 : _GEN_146; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_148 = 8'h94 == io_addr ? 8'h0 : _GEN_147; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_149 = 8'h95 == io_addr ? 8'h0 : _GEN_148; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_150 = 8'h96 == io_addr ? 8'h0 : _GEN_149; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_151 = 8'h97 == io_addr ? 8'h0 : _GEN_150; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_152 = 8'h98 == io_addr ? 8'h0 : _GEN_151; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_153 = 8'h99 == io_addr ? 8'h0 : _GEN_152; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_154 = 8'h9a == io_addr ? 8'h0 : _GEN_153; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_155 = 8'h9b == io_addr ? 8'h0 : _GEN_154; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_156 = 8'h9c == io_addr ? 8'h0 : _GEN_155; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_157 = 8'h9d == io_addr ? 8'h0 : _GEN_156; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_158 = 8'h9e == io_addr ? 8'h0 : _GEN_157; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_159 = 8'h9f == io_addr ? 8'h0 : _GEN_158; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_160 = 8'ha0 == io_addr ? 8'h0 : _GEN_159; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_161 = 8'ha1 == io_addr ? 8'h0 : _GEN_160; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_162 = 8'ha2 == io_addr ? 8'h0 : _GEN_161; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_163 = 8'ha3 == io_addr ? 8'h0 : _GEN_162; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_164 = 8'ha4 == io_addr ? 8'h0 : _GEN_163; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_165 = 8'ha5 == io_addr ? 8'h0 : _GEN_164; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_166 = 8'ha6 == io_addr ? 8'h0 : _GEN_165; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_167 = 8'ha7 == io_addr ? 8'h0 : _GEN_166; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_168 = 8'ha8 == io_addr ? 8'h0 : _GEN_167; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_169 = 8'ha9 == io_addr ? 8'h0 : _GEN_168; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_170 = 8'haa == io_addr ? 8'h0 : _GEN_169; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_171 = 8'hab == io_addr ? 8'h0 : _GEN_170; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_172 = 8'hac == io_addr ? 8'h0 : _GEN_171; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_173 = 8'had == io_addr ? 8'h0 : _GEN_172; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_174 = 8'hae == io_addr ? 8'h0 : _GEN_173; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_175 = 8'haf == io_addr ? 8'h0 : _GEN_174; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_176 = 8'hb0 == io_addr ? 8'h0 : _GEN_175; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_177 = 8'hb1 == io_addr ? 8'h0 : _GEN_176; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_178 = 8'hb2 == io_addr ? 8'h0 : _GEN_177; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_179 = 8'hb3 == io_addr ? 8'h0 : _GEN_178; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_180 = 8'hb4 == io_addr ? 8'h0 : _GEN_179; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_181 = 8'hb5 == io_addr ? 8'h0 : _GEN_180; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_182 = 8'hb6 == io_addr ? 8'h0 : _GEN_181; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_183 = 8'hb7 == io_addr ? 8'h0 : _GEN_182; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_184 = 8'hb8 == io_addr ? 8'h0 : _GEN_183; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_185 = 8'hb9 == io_addr ? 8'h0 : _GEN_184; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_186 = 8'hba == io_addr ? 8'h0 : _GEN_185; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_187 = 8'hbb == io_addr ? 8'h0 : _GEN_186; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_188 = 8'hbc == io_addr ? 8'h0 : _GEN_187; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_189 = 8'hbd == io_addr ? 8'h0 : _GEN_188; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_190 = 8'hbe == io_addr ? 8'h0 : _GEN_189; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_191 = 8'hbf == io_addr ? 8'h0 : _GEN_190; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_192 = 8'hc0 == io_addr ? 8'h0 : _GEN_191; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_193 = 8'hc1 == io_addr ? 8'h0 : _GEN_192; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_194 = 8'hc2 == io_addr ? 8'h0 : _GEN_193; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_195 = 8'hc3 == io_addr ? 8'h0 : _GEN_194; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_196 = 8'hc4 == io_addr ? 8'h0 : _GEN_195; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_197 = 8'hc5 == io_addr ? 8'h0 : _GEN_196; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_198 = 8'hc6 == io_addr ? 8'h0 : _GEN_197; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_199 = 8'hc7 == io_addr ? 8'h0 : _GEN_198; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_200 = 8'hc8 == io_addr ? 8'h0 : _GEN_199; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_201 = 8'hc9 == io_addr ? 8'h0 : _GEN_200; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_202 = 8'hca == io_addr ? 8'h0 : _GEN_201; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_203 = 8'hcb == io_addr ? 8'h0 : _GEN_202; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_204 = 8'hcc == io_addr ? 8'h0 : _GEN_203; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_205 = 8'hcd == io_addr ? 8'h0 : _GEN_204; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_206 = 8'hce == io_addr ? 8'h0 : _GEN_205; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_207 = 8'hcf == io_addr ? 8'h0 : _GEN_206; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_208 = 8'hd0 == io_addr ? 8'h0 : _GEN_207; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_209 = 8'hd1 == io_addr ? 8'h0 : _GEN_208; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_210 = 8'hd2 == io_addr ? 8'h0 : _GEN_209; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_211 = 8'hd3 == io_addr ? 8'h0 : _GEN_210; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_212 = 8'hd4 == io_addr ? 8'h0 : _GEN_211; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_213 = 8'hd5 == io_addr ? 8'h0 : _GEN_212; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_214 = 8'hd6 == io_addr ? 8'h0 : _GEN_213; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_215 = 8'hd7 == io_addr ? 8'h0 : _GEN_214; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_216 = 8'hd8 == io_addr ? 8'h0 : _GEN_215; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_217 = 8'hd9 == io_addr ? 8'h0 : _GEN_216; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_218 = 8'hda == io_addr ? 8'h0 : _GEN_217; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_219 = 8'hdb == io_addr ? 8'h0 : _GEN_218; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_220 = 8'hdc == io_addr ? 8'h0 : _GEN_219; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_221 = 8'hdd == io_addr ? 8'h0 : _GEN_220; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_222 = 8'hde == io_addr ? 8'h0 : _GEN_221; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_223 = 8'hdf == io_addr ? 8'h0 : _GEN_222; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_224 = 8'he0 == io_addr ? 8'h0 : _GEN_223; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_225 = 8'he1 == io_addr ? 8'h0 : _GEN_224; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_226 = 8'he2 == io_addr ? 8'h0 : _GEN_225; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_227 = 8'he3 == io_addr ? 8'h0 : _GEN_226; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_228 = 8'he4 == io_addr ? 8'h0 : _GEN_227; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_229 = 8'he5 == io_addr ? 8'h0 : _GEN_228; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_230 = 8'he6 == io_addr ? 8'h0 : _GEN_229; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_231 = 8'he7 == io_addr ? 8'h0 : _GEN_230; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_232 = 8'he8 == io_addr ? 8'h0 : _GEN_231; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_233 = 8'he9 == io_addr ? 8'h0 : _GEN_232; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_234 = 8'hea == io_addr ? 8'h0 : _GEN_233; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_235 = 8'heb == io_addr ? 8'h0 : _GEN_234; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_236 = 8'hec == io_addr ? 8'h0 : _GEN_235; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_237 = 8'hed == io_addr ? 8'h0 : _GEN_236; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_238 = 8'hee == io_addr ? 8'h0 : _GEN_237; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_239 = 8'hef == io_addr ? 8'h0 : _GEN_238; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_240 = 8'hf0 == io_addr ? 8'h0 : _GEN_239; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_241 = 8'hf1 == io_addr ? 8'h0 : _GEN_240; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_242 = 8'hf2 == io_addr ? 8'h0 : _GEN_241; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_243 = 8'hf3 == io_addr ? 8'h0 : _GEN_242; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_244 = 8'hf4 == io_addr ? 8'h0 : _GEN_243; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_245 = 8'hf5 == io_addr ? 8'h0 : _GEN_244; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_246 = 8'hf6 == io_addr ? 8'h0 : _GEN_245; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_247 = 8'hf7 == io_addr ? 8'h0 : _GEN_246; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_248 = 8'hf8 == io_addr ? 8'h0 : _GEN_247; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_249 = 8'hf9 == io_addr ? 8'h0 : _GEN_248; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_250 = 8'hfa == io_addr ? 8'h0 : _GEN_249; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_251 = 8'hfb == io_addr ? 8'h0 : _GEN_250; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_252 = 8'hfc == io_addr ? 8'h0 : _GEN_251; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_253 = 8'hfd == io_addr ? 8'h0 : _GEN_252; // @[Hello.scala 31:{13,13}]
  wire [7:0] _GEN_254 = 8'hfe == io_addr ? 8'h0 : _GEN_253; // @[Hello.scala 31:{13,13}]
  assign io_data = 8'hff == io_addr ? 8'h0 : _GEN_254; // @[Hello.scala 31:{13,13}]
endmodule
